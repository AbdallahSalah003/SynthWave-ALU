module carry_look_ahead_adder(
	input [31:0] A,
	input [31:0] B,
	input Cin,
	output [31:0] Sum,
	output Cout);
	wire [31:0] G, P,C;
	assign G = A & B;
	assign P = A ^ B;
	assign C[0] = G[0] | (P[0] & Cin);
	assign C[1] = G[1] | (P[1]&G[0]) | (P[1]&P[0]&Cin);
	assign C[2] = G[2] | (P[2]&G[1]) | (P[2]&P[1]&G[0]) | (P[2]&P[1]&P[0]&Cin);
	assign C[3] = G[3] | (P[3]&G[2]) | (P[3]&P[2]&G[1]) | (P[3]&P[2]&P[1]&G[0]) | (P[3]&P[2]&P[1]&P[0]&Cin);
	assign C[4] = G[4] | (P[4]&G[3]) | (P[4]&P[3]&G[2]) | (P[4]&P[3]&P[2]&G[1]) | (P[4]&P[3]&P[2]&P[1]&G[0]) | (P[4]&P[3]&P[2]&P[1]&P[0]&Cin);
	assign C[5] = G[5] | (P[5]&G[4]) | (P[5]&P[4]&G[3]) | (P[5]&P[4]&P[3]&G[2]) | (P[5]&P[4]&P[3]&P[2]&G[1]) | (P[5]&P[4]&P[3]&P[2]&P[1]&G[0]) | (P[5]&P[4]&P[3]&P[2]&P[1]&P[0]&Cin);
	assign C[6] = G[6] | (P[6]&G[5]) | (P[6]&P[5]&G[4]) | (P[6]&P[5]&P[4]&G[3]) | (P[6]&P[5]&P[4]&P[3]&G[2]) | (P[6]&P[5]&P[4]&P[3]&P[2]&G[1]) | (P[6]&P[5]&P[4]&P[3]&P[2]&P[1]&G[0]) | (P[6]&P[5]&P[4]&P[3]&P[2]&P[1]&P[0]&Cin);
	assign C[7] = G[7] | (P[7]&G[6]) | (P[7]&P[6]&G[5]) | (P[7]&P[6]&P[5]&G[4]) | (P[7]&P[6]&P[5]&P[4]&G[3]) | (P[7]&P[6]&P[5]&P[4]&P[3]&G[2]) | (P[7]&P[6]&P[5]&P[4]&P[3]&P[2]&G[1]) | (P[7]&P[6]&P[5]&P[4]&P[3]&P[2]&P[1]&G[0]) | (P[7]&P[6]&P[5]&P[4]&P[3]&P[2]&P[1]&P[0]&Cin);
	assign C[8] = G[8] | (P[8]&G[7]) | (P[8]&P[7]&G[6]) | (P[8]&P[7]&P[6]&G[5]) | (P[8]&P[7]&P[6]&P[5]&G[4]) | (P[8]&P[7]&P[6]&P[5]&P[4]&G[3]) | (P[8]&P[7]&P[6]&P[5]&P[4]&P[3]&G[2]) | (P[8]&P[7]&P[6]&P[5]&P[4]&P[3]&P[2]&G[1]) | (P[8]&P[7]&P[6]&P[5]&P[4]&P[3]&P[2]&P[1]&G[0]) | (P[8]&P[7]&P[6]&P[5]&P[4]&P[3]&P[2]&P[1]&P[0]&Cin);
	assign C[9] = G[9] | (P[9]&G[8]) | (P[9]&P[8]&G[7]) | (P[9]&P[8]&P[7]&G[6]) | (P[9]&P[8]&P[7]&P[6]&G[5]) | (P[9]&P[8]&P[7]&P[6]&P[5]&G[4]) | (P[9]&P[8]&P[7]&P[6]&P[5]&P[4]&G[3]) | (P[9]&P[8]&P[7]&P[6]&P[5]&P[4]&P[3]&G[2]) | (P[9]&P[8]&P[7]&P[6]&P[5]&P[4]&P[3]&P[2]&G[1]) | (P[9]&P[8]&P[7]&P[6]&P[5]&P[4]&P[3]&P[2]&P[1]&G[0]) | (P[9]&P[8]&P[7]&P[6]&P[5]&P[4]&P[3]&P[2]&P[1]&P[0]&Cin);
	assign C[10] = G[10] | (P[10]&G[9]) | (P[10]&P[9]&G[8]) | (P[10]&P[9]&P[8]&G[7]) | (P[10]&P[9]&P[8]&P[7]&G[6]) | (P[10]&P[9]&P[8]&P[7]&P[6]&G[5]) | (P[10]&P[9]&P[8]&P[7]&P[6]&P[5]&G[4]) | (P[10]&P[9]&P[8]&P[7]&P[6]&P[5]&P[4]&G[3]) | (P[10]&P[9]&P[8]&P[7]&P[6]&P[5]&P[4]&P[3]&G[2]) | (P[10]&P[9]&P[8]&P[7]&P[6]&P[5]&P[4]&P[3]&P[2]&G[1]) | (P[10]&P[9]&P[8]&P[7]&P[6]&P[5]&P[4]&P[3]&P[2]&P[1]&G[0]) | (P[10]&P[9]&P[8]&P[7]&P[6]&P[5]&P[4]&P[3]&P[2]&P[1]&P[0]&Cin);
	assign C[11] = G[11] | (P[11]&G[10]) | (P[11]&P[10]&G[9]) | (P[11]&P[10]&P[9]&G[8]) | (P[11]&P[10]&P[9]&P[8]&G[7]) | (P[11]&P[10]&P[9]&P[8]&P[7]&G[6]) | (P[11]&P[10]&P[9]&P[8]&P[7]&P[6]&G[5]) | (P[11]&P[10]&P[9]&P[8]&P[7]&P[6]&P[5]&G[4]) | (P[11]&P[10]&P[9]&P[8]&P[7]&P[6]&P[5]&P[4]&G[3]) | (P[11]&P[10]&P[9]&P[8]&P[7]&P[6]&P[5]&P[4]&P[3]&G[2]) | (P[11]&P[10]&P[9]&P[8]&P[7]&P[6]&P[5]&P[4]&P[3]&P[2]&G[1]) | (P[11]&P[10]&P[9]&P[8]&P[7]&P[6]&P[5]&P[4]&P[3]&P[2]&P[1]&G[0]) | (P[11]&P[10]&P[9]&P[8]&P[7]&P[6]&P[5]&P[4]&P[3]&P[2]&P[1]&P[0]&Cin);
	assign C[12] = G[12] | (P[12]&G[11]) | (P[12]&P[11]&G[10]) | (P[12]&P[11]&P[10]&G[9]) | (P[12]&P[11]&P[10]&P[9]&G[8]) | (P[12]&P[11]&P[10]&P[9]&P[8]&G[7]) | (P[12]&P[11]&P[10]&P[9]&P[8]&P[7]&G[6]) | (P[12]&P[11]&P[10]&P[9]&P[8]&P[7]&P[6]&G[5]) | (P[12]&P[11]&P[10]&P[9]&P[8]&P[7]&P[6]&P[5]&G[4]) | (P[12]&P[11]&P[10]&P[9]&P[8]&P[7]&P[6]&P[5]&P[4]&G[3]) | (P[12]&P[11]&P[10]&P[9]&P[8]&P[7]&P[6]&P[5]&P[4]&P[3]&G[2]) | (P[12]&P[11]&P[10]&P[9]&P[8]&P[7]&P[6]&P[5]&P[4]&P[3]&P[2]&G[1]) | (P[12]&P[11]&P[10]&P[9]&P[8]&P[7]&P[6]&P[5]&P[4]&P[3]&P[2]&P[1]&G[0]) | (P[12]&P[11]&P[10]&P[9]&P[8]&P[7]&P[6]&P[5]&P[4]&P[3]&P[2]&P[1]&P[0]&Cin);
	assign C[13] = G[13] | (P[13]&G[12]) | (P[13]&P[12]&G[11]) | (P[13]&P[12]&P[11]&G[10]) | (P[13]&P[12]&P[11]&P[10]&G[9]) | (P[13]&P[12]&P[11]&P[10]&P[9]&G[8]) | (P[13]&P[12]&P[11]&P[10]&P[9]&P[8]&G[7]) | (P[13]&P[12]&P[11]&P[10]&P[9]&P[8]&P[7]&G[6]) | (P[13]&P[12]&P[11]&P[10]&P[9]&P[8]&P[7]&P[6]&G[5]) | (P[13]&P[12]&P[11]&P[10]&P[9]&P[8]&P[7]&P[6]&P[5]&G[4]) | (P[13]&P[12]&P[11]&P[10]&P[9]&P[8]&P[7]&P[6]&P[5]&P[4]&G[3]) | (P[13]&P[12]&P[11]&P[10]&P[9]&P[8]&P[7]&P[6]&P[5]&P[4]&P[3]&G[2]) | (P[13]&P[12]&P[11]&P[10]&P[9]&P[8]&P[7]&P[6]&P[5]&P[4]&P[3]&P[2]&G[1]) | (P[13]&P[12]&P[11]&P[10]&P[9]&P[8]&P[7]&P[6]&P[5]&P[4]&P[3]&P[2]&P[1]&G[0]) | (P[13]&P[12]&P[11]&P[10]&P[9]&P[8]&P[7]&P[6]&P[5]&P[4]&P[3]&P[2]&P[1]&P[0]&Cin);
	assign C[14] = G[14] | (P[14]&G[13]) | (P[14]&P[13]&G[12]) | (P[14]&P[13]&P[12]&G[11]) | (P[14]&P[13]&P[12]&P[11]&G[10]) | (P[14]&P[13]&P[12]&P[11]&P[10]&G[9]) | (P[14]&P[13]&P[12]&P[11]&P[10]&P[9]&G[8]) | (P[14]&P[13]&P[12]&P[11]&P[10]&P[9]&P[8]&G[7]) | (P[14]&P[13]&P[12]&P[11]&P[10]&P[9]&P[8]&P[7]&G[6]) | (P[14]&P[13]&P[12]&P[11]&P[10]&P[9]&P[8]&P[7]&P[6]&G[5]) | (P[14]&P[13]&P[12]&P[11]&P[10]&P[9]&P[8]&P[7]&P[6]&P[5]&G[4]) | (P[14]&P[13]&P[12]&P[11]&P[10]&P[9]&P[8]&P[7]&P[6]&P[5]&P[4]&G[3]) | (P[14]&P[13]&P[12]&P[11]&P[10]&P[9]&P[8]&P[7]&P[6]&P[5]&P[4]&P[3]&G[2]) | (P[14]&P[13]&P[12]&P[11]&P[10]&P[9]&P[8]&P[7]&P[6]&P[5]&P[4]&P[3]&P[2]&G[1]) | (P[14]&P[13]&P[12]&P[11]&P[10]&P[9]&P[8]&P[7]&P[6]&P[5]&P[4]&P[3]&P[2]&P[1]&G[0]) | (P[14]&P[13]&P[12]&P[11]&P[10]&P[9]&P[8]&P[7]&P[6]&P[5]&P[4]&P[3]&P[2]&P[1]&P[0]&Cin);
	assign C[15] = G[15] | (P[15]&G[14]) | (P[15]&P[14]&G[13]) | (P[15]&P[14]&P[13]&G[12]) | (P[15]&P[14]&P[13]&P[12]&G[11]) | (P[15]&P[14]&P[13]&P[12]&P[11]&G[10]) | (P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&G[9]) | (P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&P[9]&G[8]) | (P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&P[9]&P[8]&G[7]) | (P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&P[9]&P[8]&P[7]&G[6]) | (P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&P[9]&P[8]&P[7]&P[6]&G[5]) | (P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&P[9]&P[8]&P[7]&P[6]&P[5]&G[4]) | (P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&P[9]&P[8]&P[7]&P[6]&P[5]&P[4]&G[3]) | (P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&P[9]&P[8]&P[7]&P[6]&P[5]&P[4]&P[3]&G[2]) | (P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&P[9]&P[8]&P[7]&P[6]&P[5]&P[4]&P[3]&P[2]&G[1]) | (P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&P[9]&P[8]&P[7]&P[6]&P[5]&P[4]&P[3]&P[2]&P[1]&G[0]) | (P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&P[9]&P[8]&P[7]&P[6]&P[5]&P[4]&P[3]&P[2]&P[1]&P[0]&Cin);
	assign C[16] = G[16] | (P[16]&G[15]) | (P[16]&P[15]&G[14]) | (P[16]&P[15]&P[14]&G[13]) | (P[16]&P[15]&P[14]&P[13]&G[12]) | (P[16]&P[15]&P[14]&P[13]&P[12]&G[11]) | (P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&G[10]) | (P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&G[9]) | (P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&P[9]&G[8]) | (P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&P[9]&P[8]&G[7]) | (P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&P[9]&P[8]&P[7]&G[6]) | (P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&P[9]&P[8]&P[7]&P[6]&G[5]) | (P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&P[9]&P[8]&P[7]&P[6]&P[5]&G[4]) | (P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&P[9]&P[8]&P[7]&P[6]&P[5]&P[4]&G[3]) | (P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&P[9]&P[8]&P[7]&P[6]&P[5]&P[4]&P[3]&G[2]) | (P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&P[9]&P[8]&P[7]&P[6]&P[5]&P[4]&P[3]&P[2]&G[1]) | (P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&P[9]&P[8]&P[7]&P[6]&P[5]&P[4]&P[3]&P[2]&P[1]&G[0]) | (P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&P[9]&P[8]&P[7]&P[6]&P[5]&P[4]&P[3]&P[2]&P[1]&P[0]&Cin);
	assign C[17] = G[17] | (P[17]&G[16]) | (P[17]&P[16]&G[15]) | (P[17]&P[16]&P[15]&G[14]) | (P[17]&P[16]&P[15]&P[14]&G[13]) | (P[17]&P[16]&P[15]&P[14]&P[13]&G[12]) | (P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&G[11]) | (P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&G[10]) | (P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&G[9]) | (P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&P[9]&G[8]) | (P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&P[9]&P[8]&G[7]) | (P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&P[9]&P[8]&P[7]&G[6]) | (P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&P[9]&P[8]&P[7]&P[6]&G[5]) | (P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&P[9]&P[8]&P[7]&P[6]&P[5]&G[4]) | (P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&P[9]&P[8]&P[7]&P[6]&P[5]&P[4]&G[3]) | (P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&P[9]&P[8]&P[7]&P[6]&P[5]&P[4]&P[3]&G[2]) | (P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&P[9]&P[8]&P[7]&P[6]&P[5]&P[4]&P[3]&P[2]&G[1]) | (P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&P[9]&P[8]&P[7]&P[6]&P[5]&P[4]&P[3]&P[2]&P[1]&G[0]) | (P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&P[9]&P[8]&P[7]&P[6]&P[5]&P[4]&P[3]&P[2]&P[1]&P[0]&Cin);
	assign C[18] = G[18] | (P[18]&G[17]) | (P[18]&P[17]&G[16]) | (P[18]&P[17]&P[16]&G[15]) | (P[18]&P[17]&P[16]&P[15]&G[14]) | (P[18]&P[17]&P[16]&P[15]&P[14]&G[13]) | (P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&G[12]) | (P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&G[11]) | (P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&G[10]) | (P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&G[9]) | (P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&P[9]&G[8]) | (P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&P[9]&P[8]&G[7]) | (P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&P[9]&P[8]&P[7]&G[6]) | (P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&P[9]&P[8]&P[7]&P[6]&G[5]) | (P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&P[9]&P[8]&P[7]&P[6]&P[5]&G[4]) | (P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&P[9]&P[8]&P[7]&P[6]&P[5]&P[4]&G[3]) | (P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&P[9]&P[8]&P[7]&P[6]&P[5]&P[4]&P[3]&G[2]) | (P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&P[9]&P[8]&P[7]&P[6]&P[5]&P[4]&P[3]&P[2]&G[1]) | (P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&P[9]&P[8]&P[7]&P[6]&P[5]&P[4]&P[3]&P[2]&P[1]&G[0]) | (P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&P[9]&P[8]&P[7]&P[6]&P[5]&P[4]&P[3]&P[2]&P[1]&P[0]&Cin);
	assign C[19] = G[19] | (P[19]&G[18]) | (P[19]&P[18]&G[17]) | (P[19]&P[18]&P[17]&G[16]) | (P[19]&P[18]&P[17]&P[16]&G[15]) | (P[19]&P[18]&P[17]&P[16]&P[15]&G[14]) | (P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&G[13]) | (P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&G[12]) | (P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&G[11]) | (P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&G[10]) | (P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&G[9]) | (P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&P[9]&G[8]) | (P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&P[9]&P[8]&G[7]) | (P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&P[9]&P[8]&P[7]&G[6]) | (P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&P[9]&P[8]&P[7]&P[6]&G[5]) | (P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&P[9]&P[8]&P[7]&P[6]&P[5]&G[4]) | (P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&P[9]&P[8]&P[7]&P[6]&P[5]&P[4]&G[3]) | (P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&P[9]&P[8]&P[7]&P[6]&P[5]&P[4]&P[3]&G[2]) | (P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&P[9]&P[8]&P[7]&P[6]&P[5]&P[4]&P[3]&P[2]&G[1]) | (P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&P[9]&P[8]&P[7]&P[6]&P[5]&P[4]&P[3]&P[2]&P[1]&G[0]) | (P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&P[9]&P[8]&P[7]&P[6]&P[5]&P[4]&P[3]&P[2]&P[1]&P[0]&Cin);
	assign C[20] = G[20] | (P[20]&G[19]) | (P[20]&P[19]&G[18]) | (P[20]&P[19]&P[18]&G[17]) | (P[20]&P[19]&P[18]&P[17]&G[16]) | (P[20]&P[19]&P[18]&P[17]&P[16]&G[15]) | (P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&G[14]) | (P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&G[13]) | (P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&G[12]) | (P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&G[11]) | (P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&G[10]) | (P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&G[9]) | (P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&P[9]&G[8]) | (P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&P[9]&P[8]&G[7]) | (P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&P[9]&P[8]&P[7]&G[6]) | (P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&P[9]&P[8]&P[7]&P[6]&G[5]) | (P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&P[9]&P[8]&P[7]&P[6]&P[5]&G[4]) | (P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&P[9]&P[8]&P[7]&P[6]&P[5]&P[4]&G[3]) | (P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&P[9]&P[8]&P[7]&P[6]&P[5]&P[4]&P[3]&G[2]) | (P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&P[9]&P[8]&P[7]&P[6]&P[5]&P[4]&P[3]&P[2]&G[1]) | (P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&P[9]&P[8]&P[7]&P[6]&P[5]&P[4]&P[3]&P[2]&P[1]&G[0]) | (P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&P[9]&P[8]&P[7]&P[6]&P[5]&P[4]&P[3]&P[2]&P[1]&P[0]&Cin);
	assign C[21] = G[21] | (P[21]&G[20]) | (P[21]&P[20]&G[19]) | (P[21]&P[20]&P[19]&G[18]) | (P[21]&P[20]&P[19]&P[18]&G[17]) | (P[21]&P[20]&P[19]&P[18]&P[17]&G[16]) | (P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&G[15]) | (P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&G[14]) | (P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&G[13]) | (P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&G[12]) | (P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&G[11]) | (P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&G[10]) | (P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&G[9]) | (P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&P[9]&G[8]) | (P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&P[9]&P[8]&G[7]) | (P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&P[9]&P[8]&P[7]&G[6]) | (P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&P[9]&P[8]&P[7]&P[6]&G[5]) | (P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&P[9]&P[8]&P[7]&P[6]&P[5]&G[4]) | (P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&P[9]&P[8]&P[7]&P[6]&P[5]&P[4]&G[3]) | (P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&P[9]&P[8]&P[7]&P[6]&P[5]&P[4]&P[3]&G[2]) | (P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&P[9]&P[8]&P[7]&P[6]&P[5]&P[4]&P[3]&P[2]&G[1]) | (P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&P[9]&P[8]&P[7]&P[6]&P[5]&P[4]&P[3]&P[2]&P[1]&G[0]) | (P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&P[9]&P[8]&P[7]&P[6]&P[5]&P[4]&P[3]&P[2]&P[1]&P[0]&Cin);
	assign C[22] = G[22] | (P[22]&G[21]) | (P[22]&P[21]&G[20]) | (P[22]&P[21]&P[20]&G[19]) | (P[22]&P[21]&P[20]&P[19]&G[18]) | (P[22]&P[21]&P[20]&P[19]&P[18]&G[17]) | (P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&G[16]) | (P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&G[15]) | (P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&G[14]) | (P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&G[13]) | (P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&G[12]) | (P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&G[11]) | (P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&G[10]) | (P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&G[9]) | (P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&P[9]&G[8]) | (P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&P[9]&P[8]&G[7]) | (P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&P[9]&P[8]&P[7]&G[6]) | (P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&P[9]&P[8]&P[7]&P[6]&G[5]) | (P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&P[9]&P[8]&P[7]&P[6]&P[5]&G[4]) | (P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&P[9]&P[8]&P[7]&P[6]&P[5]&P[4]&G[3]) | (P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&P[9]&P[8]&P[7]&P[6]&P[5]&P[4]&P[3]&G[2]) | (P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&P[9]&P[8]&P[7]&P[6]&P[5]&P[4]&P[3]&P[2]&G[1]) | (P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&P[9]&P[8]&P[7]&P[6]&P[5]&P[4]&P[3]&P[2]&P[1]&G[0]) | (P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&P[9]&P[8]&P[7]&P[6]&P[5]&P[4]&P[3]&P[2]&P[1]&P[0]&Cin);
	assign C[23] = G[23] | (P[23]&G[22]) | (P[23]&P[22]&G[21]) | (P[23]&P[22]&P[21]&G[20]) | (P[23]&P[22]&P[21]&P[20]&G[19]) | (P[23]&P[22]&P[21]&P[20]&P[19]&G[18]) | (P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&G[17]) | (P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&G[16]) | (P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&G[15]) | (P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&G[14]) | (P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&G[13]) | (P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&G[12]) | (P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&G[11]) | (P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&G[10]) | (P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&G[9]) | (P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&P[9]&G[8]) | (P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&P[9]&P[8]&G[7]) | (P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&P[9]&P[8]&P[7]&G[6]) | (P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&P[9]&P[8]&P[7]&P[6]&G[5]) | (P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&P[9]&P[8]&P[7]&P[6]&P[5]&G[4]) | (P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&P[9]&P[8]&P[7]&P[6]&P[5]&P[4]&G[3]) | (P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&P[9]&P[8]&P[7]&P[6]&P[5]&P[4]&P[3]&G[2]) | (P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&P[9]&P[8]&P[7]&P[6]&P[5]&P[4]&P[3]&P[2]&G[1]) | (P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&P[9]&P[8]&P[7]&P[6]&P[5]&P[4]&P[3]&P[2]&P[1]&G[0]) | (P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&P[9]&P[8]&P[7]&P[6]&P[5]&P[4]&P[3]&P[2]&P[1]&P[0]&Cin);
	assign C[24] = G[24] | (P[24]&G[23]) | (P[24]&P[23]&G[22]) | (P[24]&P[23]&P[22]&G[21]) | (P[24]&P[23]&P[22]&P[21]&G[20]) | (P[24]&P[23]&P[22]&P[21]&P[20]&G[19]) | (P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&G[18]) | (P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&G[17]) | (P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&G[16]) | (P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&G[15]) | (P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&G[14]) | (P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&G[13]) | (P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&G[12]) | (P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&G[11]) | (P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&G[10]) | (P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&G[9]) | (P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&P[9]&G[8]) | (P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&P[9]&P[8]&G[7]) | (P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&P[9]&P[8]&P[7]&G[6]) | (P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&P[9]&P[8]&P[7]&P[6]&G[5]) | (P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&P[9]&P[8]&P[7]&P[6]&P[5]&G[4]) | (P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&P[9]&P[8]&P[7]&P[6]&P[5]&P[4]&G[3]) | (P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&P[9]&P[8]&P[7]&P[6]&P[5]&P[4]&P[3]&G[2]) | (P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&P[9]&P[8]&P[7]&P[6]&P[5]&P[4]&P[3]&P[2]&G[1]) | (P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&P[9]&P[8]&P[7]&P[6]&P[5]&P[4]&P[3]&P[2]&P[1]&G[0]) | (P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&P[9]&P[8]&P[7]&P[6]&P[5]&P[4]&P[3]&P[2]&P[1]&P[0]&Cin);
	assign C[25] = G[25] | (P[25]&G[24]) | (P[25]&P[24]&G[23]) | (P[25]&P[24]&P[23]&G[22]) | (P[25]&P[24]&P[23]&P[22]&G[21]) | (P[25]&P[24]&P[23]&P[22]&P[21]&G[20]) | (P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&G[19]) | (P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&G[18]) | (P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&G[17]) | (P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&G[16]) | (P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&G[15]) | (P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&G[14]) | (P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&G[13]) | (P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&G[12]) | (P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&G[11]) | (P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&G[10]) | (P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&G[9]) | (P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&P[9]&G[8]) | (P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&P[9]&P[8]&G[7]) | (P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&P[9]&P[8]&P[7]&G[6]) | (P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&P[9]&P[8]&P[7]&P[6]&G[5]) | (P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&P[9]&P[8]&P[7]&P[6]&P[5]&G[4]) | (P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&P[9]&P[8]&P[7]&P[6]&P[5]&P[4]&G[3]) | (P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&P[9]&P[8]&P[7]&P[6]&P[5]&P[4]&P[3]&G[2]) | (P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&P[9]&P[8]&P[7]&P[6]&P[5]&P[4]&P[3]&P[2]&G[1]) | (P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&P[9]&P[8]&P[7]&P[6]&P[5]&P[4]&P[3]&P[2]&P[1]&G[0]) | (P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&P[9]&P[8]&P[7]&P[6]&P[5]&P[4]&P[3]&P[2]&P[1]&P[0]&Cin);
	assign C[26] = G[26] | (P[26]&G[25]) | (P[26]&P[25]&G[24]) | (P[26]&P[25]&P[24]&G[23]) | (P[26]&P[25]&P[24]&P[23]&G[22]) | (P[26]&P[25]&P[24]&P[23]&P[22]&G[21]) | (P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&G[20]) | (P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&G[19]) | (P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&G[18]) | (P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&G[17]) | (P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&G[16]) | (P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&G[15]) | (P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&G[14]) | (P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&G[13]) | (P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&G[12]) | (P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&G[11]) | (P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&G[10]) | (P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&G[9]) | (P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&P[9]&G[8]) | (P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&P[9]&P[8]&G[7]) | (P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&P[9]&P[8]&P[7]&G[6]) | (P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&P[9]&P[8]&P[7]&P[6]&G[5]) | (P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&P[9]&P[8]&P[7]&P[6]&P[5]&G[4]) | (P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&P[9]&P[8]&P[7]&P[6]&P[5]&P[4]&G[3]) | (P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&P[9]&P[8]&P[7]&P[6]&P[5]&P[4]&P[3]&G[2]) | (P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&P[9]&P[8]&P[7]&P[6]&P[5]&P[4]&P[3]&P[2]&G[1]) | (P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&P[9]&P[8]&P[7]&P[6]&P[5]&P[4]&P[3]&P[2]&P[1]&G[0]) | (P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&P[9]&P[8]&P[7]&P[6]&P[5]&P[4]&P[3]&P[2]&P[1]&P[0]&Cin);
	assign C[27] = G[27] | (P[27]&G[26]) | (P[27]&P[26]&G[25]) | (P[27]&P[26]&P[25]&G[24]) | (P[27]&P[26]&P[25]&P[24]&G[23]) | (P[27]&P[26]&P[25]&P[24]&P[23]&G[22]) | (P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&G[21]) | (P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&G[20]) | (P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&G[19]) | (P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&G[18]) | (P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&G[17]) | (P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&G[16]) | (P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&G[15]) | (P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&G[14]) | (P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&G[13]) | (P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&G[12]) | (P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&G[11]) | (P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&G[10]) | (P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&G[9]) | (P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&P[9]&G[8]) | (P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&P[9]&P[8]&G[7]) | (P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&P[9]&P[8]&P[7]&G[6]) | (P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&P[9]&P[8]&P[7]&P[6]&G[5]) | (P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&P[9]&P[8]&P[7]&P[6]&P[5]&G[4]) | (P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&P[9]&P[8]&P[7]&P[6]&P[5]&P[4]&G[3]) | (P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&P[9]&P[8]&P[7]&P[6]&P[5]&P[4]&P[3]&G[2]) | (P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&P[9]&P[8]&P[7]&P[6]&P[5]&P[4]&P[3]&P[2]&G[1]) | (P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&P[9]&P[8]&P[7]&P[6]&P[5]&P[4]&P[3]&P[2]&P[1]&G[0]) | (P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&P[9]&P[8]&P[7]&P[6]&P[5]&P[4]&P[3]&P[2]&P[1]&P[0]&Cin);
	assign C[28] = G[28] | (P[28]&G[27]) | (P[28]&P[27]&G[26]) | (P[28]&P[27]&P[26]&G[25]) | (P[28]&P[27]&P[26]&P[25]&G[24]) | (P[28]&P[27]&P[26]&P[25]&P[24]&G[23]) | (P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&G[22]) | (P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&G[21]) | (P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&G[20]) | (P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&G[19]) | (P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&G[18]) | (P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&G[17]) | (P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&G[16]) | (P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&G[15]) | (P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&G[14]) | (P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&G[13]) | (P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&G[12]) | (P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&G[11]) | (P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&G[10]) | (P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&G[9]) | (P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&P[9]&G[8]) | (P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&P[9]&P[8]&G[7]) | (P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&P[9]&P[8]&P[7]&G[6]) | (P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&P[9]&P[8]&P[7]&P[6]&G[5]) | (P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&P[9]&P[8]&P[7]&P[6]&P[5]&G[4]) | (P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&P[9]&P[8]&P[7]&P[6]&P[5]&P[4]&G[3]) | (P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&P[9]&P[8]&P[7]&P[6]&P[5]&P[4]&P[3]&G[2]) | (P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&P[9]&P[8]&P[7]&P[6]&P[5]&P[4]&P[3]&P[2]&G[1]) | (P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&P[9]&P[8]&P[7]&P[6]&P[5]&P[4]&P[3]&P[2]&P[1]&G[0]) | (P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&P[9]&P[8]&P[7]&P[6]&P[5]&P[4]&P[3]&P[2]&P[1]&P[0]&Cin);
	assign C[29] = G[29] | (P[29]&G[28]) | (P[29]&P[28]&G[27]) | (P[29]&P[28]&P[27]&G[26]) | (P[29]&P[28]&P[27]&P[26]&G[25]) | (P[29]&P[28]&P[27]&P[26]&P[25]&G[24]) | (P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&G[23]) | (P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&G[22]) | (P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&G[21]) | (P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&G[20]) | (P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&G[19]) | (P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&G[18]) | (P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&G[17]) | (P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&G[16]) | (P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&G[15]) | (P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&G[14]) | (P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&G[13]) | (P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&G[12]) | (P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&G[11]) | (P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&G[10]) | (P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&G[9]) | (P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&P[9]&G[8]) | (P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&P[9]&P[8]&G[7]) | (P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&P[9]&P[8]&P[7]&G[6]) | (P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&P[9]&P[8]&P[7]&P[6]&G[5]) | (P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&P[9]&P[8]&P[7]&P[6]&P[5]&G[4]) | (P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&P[9]&P[8]&P[7]&P[6]&P[5]&P[4]&G[3]) | (P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&P[9]&P[8]&P[7]&P[6]&P[5]&P[4]&P[3]&G[2]) | (P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&P[9]&P[8]&P[7]&P[6]&P[5]&P[4]&P[3]&P[2]&G[1]) | (P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&P[9]&P[8]&P[7]&P[6]&P[5]&P[4]&P[3]&P[2]&P[1]&G[0]) | (P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&P[9]&P[8]&P[7]&P[6]&P[5]&P[4]&P[3]&P[2]&P[1]&P[0]&Cin);
	assign C[30] = G[30] | (P[30]&G[29]) | (P[30]&P[29]&G[28]) | (P[30]&P[29]&P[28]&G[27]) | (P[30]&P[29]&P[28]&P[27]&G[26]) | (P[30]&P[29]&P[28]&P[27]&P[26]&G[25]) | (P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&G[24]) | (P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&G[23]) | (P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&G[22]) | (P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&G[21]) | (P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&G[20]) | (P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&G[19]) | (P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&G[18]) | (P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&G[17]) | (P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&G[16]) | (P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&G[15]) | (P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&G[14]) | (P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&G[13]) | (P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&G[12]) | (P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&G[11]) | (P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&G[10]) | (P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&G[9]) | (P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&P[9]&G[8]) | (P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&P[9]&P[8]&G[7]) | (P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&P[9]&P[8]&P[7]&G[6]) | (P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&P[9]&P[8]&P[7]&P[6]&G[5]) | (P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&P[9]&P[8]&P[7]&P[6]&P[5]&G[4]) | (P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&P[9]&P[8]&P[7]&P[6]&P[5]&P[4]&G[3]) | (P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&P[9]&P[8]&P[7]&P[6]&P[5]&P[4]&P[3]&G[2]) | (P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&P[9]&P[8]&P[7]&P[6]&P[5]&P[4]&P[3]&P[2]&G[1]) | (P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&P[9]&P[8]&P[7]&P[6]&P[5]&P[4]&P[3]&P[2]&P[1]&G[0]) | (P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&P[9]&P[8]&P[7]&P[6]&P[5]&P[4]&P[3]&P[2]&P[1]&P[0]&Cin);
	assign C[31] = G[31] | (P[31]&G[30]) | (P[31]&P[30]&G[29]) | (P[31]&P[30]&P[29]&G[28]) | (P[31]&P[30]&P[29]&P[28]&G[27]) | (P[31]&P[30]&P[29]&P[28]&P[27]&G[26]) | (P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&G[25]) | (P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&G[24]) | (P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&G[23]) | (P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&G[22]) | (P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&G[21]) | (P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&G[20]) | (P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&G[19]) | (P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&G[18]) | (P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&G[17]) | (P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&G[16]) | (P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&G[15]) | (P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&G[14]) | (P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&G[13]) | (P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&G[12]) | (P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&G[11]) | (P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&G[10]) | (P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&G[9]) | (P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&P[9]&G[8]) | (P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&P[9]&P[8]&G[7]) | (P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&P[9]&P[8]&P[7]&G[6]) | (P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&P[9]&P[8]&P[7]&P[6]&G[5]) | (P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&P[9]&P[8]&P[7]&P[6]&P[5]&G[4]) | (P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&P[9]&P[8]&P[7]&P[6]&P[5]&P[4]&G[3]) | (P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&P[9]&P[8]&P[7]&P[6]&P[5]&P[4]&P[3]&G[2]) | (P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&P[9]&P[8]&P[7]&P[6]&P[5]&P[4]&P[3]&P[2]&G[1]) | (P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&P[9]&P[8]&P[7]&P[6]&P[5]&P[4]&P[3]&P[2]&P[1]&G[0]) | (P[31]&P[30]&P[29]&P[28]&P[27]&P[26]&P[25]&P[24]&P[23]&P[22]&P[21]&P[20]&P[19]&P[18]&P[17]&P[16]&P[15]&P[14]&P[13]&P[12]&P[11]&P[10]&P[9]&P[8]&P[7]&P[6]&P[5]&P[4]&P[3]&P[2]&P[1]&P[0]&Cin);
	assign Sum = A ^ B ^ {C[30:0], Cin};
	assign Cout = C[31];
endmodule